
`default_nettype none
`timescale 1ns / 100ps

module tb ();

    initial begin
        $dumpfile("dsp.vcd");
        $dumpvars(0, tb);
        #500000 $finish;
    end

    reg ck = 0;

    always #42 ck <= !ck;

    reg [0:0] reset_cnt = 0;
    wire rst = & reset_cnt;

    always @(posedge ck) begin
        if (!rst)
            reset_cnt <= reset_cnt + 1;
    end

    reg        iomem_valid;
    wire       iomem_ready;
    reg [3:0]  iomem_wstrb;
    reg [31:0] iomem_addr;
    reg [31:0] iomem_wdata;
    wire [31:0] iomem_rdata;

    // Write audio test data into memory

    task write(input [31:0] addr, input [31:0] data);
        begin
            @(posedge ck);
            iomem_addr <= addr;
            iomem_wdata <= data;
            iomem_wstrb <= 4'b1111;
            iomem_valid <= 1;
            @(posedge ck);
            @(posedge ck);
        end
    endtask

    task read(input [31:0] addr);

            @(posedge ck);
            iomem_addr <= addr;
            iomem_wstrb <= 0;
            iomem_valid <= 1;
            @(posedge ck);
            @(posedge ck);

    endtask

    // Simulate removing iomem_valid
    always @(posedge ck) begin
        if (iomem_ready || !rst) begin
            iomem_valid <= 0;
            iomem_wstrb <= 0;            
            iomem_addr <= 32'hZ;
            iomem_wdata <= 32'hZ;
        end
    end

    task write_opcode;
        
        input [31:0] addr;
        input [6:0] opcode;
        input [4:0] offset;
        input [3:0] chan;
        input [15:0] gain;

        integer i;

        begin
            i = gain + (chan << 16) + (offset << 20) + (opcode << 25); 
            write(addr, i);
            $display("%h", i);
        end

    endtask

    task capture;

        input [31:0] addr;
        input [2:0] code;

        begin
            write_opcode(addr, 7'b0010000 + code, 0, 0, 0);
        end

    endtask

    task noop;

        input [31:0] addr;

        begin
            write_opcode(addr, 7'b0000000, 0, 0, 0);
        end

    endtask

    task save;

        input [31:0] addr;
        input [5:0] shift;
        input [5:0] offset;

        begin
            write_opcode(addr, 7'b1010000, 0, 0, 0);
        end

    endtask

    integer i;

    initial begin
        @(posedge ck);
        @(posedge ck);
        @(posedge ck);
        @(posedge ck);
        @(posedge ck);
        // Setup the coefficient RAM
        i = 32'h60000000;

        write(i, 32'h48000004); i += 4;
        write(i, 32'h40010004); i += 4;
        write(i, 32'h10180000); i += 4;
        write(i, 32'h48010008); i += 4;
        write(i, 32'h50000008); i += 4;
        write(i, 32'h10200001); i += 4;
        write(i, 32'h78000000); i += 4;
        write(i, 32'h78000000); i += 4;

        i = 32'h60000000;
        read(i);
 
        // set control register
        write(32'h62000000, 1); // allow_audio_writes

        // Write to audio RAM
        i = 32'h64000000;
        write(i + 0, 32'h00001234);
        write(i + 4, 32'h0000abcd);
        write(i + 8, 32'h00002323);
        write(i + (30'h40 << 2), 32'h00002222);

        write(i + (30'h44 << 2), 32'h00001111);
        write(i + (30'h45 << 2), 32'h00001234);
        write(i + (30'h46 << 2), 32'h0000abcd);
        write(i + (30'h47 << 2), 32'h00002222);

        reset_cnt <= 0;

        for (int i = 0; i < 200; i += 1) begin
            @(posedge ck);
        end
        write(32'h62000000, 0); // disable allow_audio_writes
        
    end

    /* verilator lint_off UNUSED */
    wire [7:0] test;
    /* verilator lint_on UNUSED */

    // Sync to the sck/ws I2S signals generated by the engine.
    wire sd_out, sck, ws;
    wire [5:0] frame_posn;
    wire sen;
    i2s_secondary i2sx (.ck(ck), .sck(sck), .ws(ws), .en(sen), .frame_posn(frame_posn));

    reg [15:0] left  = 16'h1234;
    reg [15:0] right = 16'habcd;

    wire sd_gen;
    i2s_tx txx(.ck(ck), .en(sen), .frame_posn(frame_posn), .sd(sd_gen), .left(left), .right(right));

    audio_engine engine(.ck(ck), .rst(rst),
        .iomem_valid(iomem_valid),
        .iomem_ready(iomem_ready),
        .iomem_wstrb(iomem_wstrb),
        .iomem_addr(iomem_addr),
        .iomem_wdata(iomem_wdata),
        .iomem_rdata(iomem_rdata),
        .sck(sck), .ws(ws),
        .sd_out(sd_out), .sd_in0(sd_gen),
        .test(test)
    );


endmodule

